library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Decodificador is
	port(
		B0, B1, B2, B3: in std_logic;
		A, B, C, D, E, F, G : out std_logic
	);
end Decodificador;

Architecture comportamento of Decodificador is
begin
	 A <= (NOT B0 AND NOT B1 AND NOT B2 AND B3) OR (NOT B0 AND B1 AND NOT B2 AND NOT B3) OR (B0 AND B1 AND NOT B2 AND B3) OR (B0 AND NOT B1 AND B2 AND B3);  
    B <= (B0 AND B2 AND B3) OR (B1 AND B2 AND NOT B3) OR (B0 AND B1 AND NOT B3) OR (NOT B0 AND B1 AND NOT B2 AND B3);
    C <= (B0 AND B1 AND B2) OR (B0 AND B1 AND NOT B3) OR (NOT B0 AND NOT B1 AND B2 AND NOT B3);
    D <= (B1 AND B2 AND B3) OR (NOT B0 AND NOT B1 AND NOT B2 AND B3) OR (NOT B0 AND B1 AND NOT B2 AND NOT B3) OR (B0 AND NOT B1 AND B2 AND NOT B3);
    E <= (NOT B0 AND B3) OR (NOT B1 AND NOT B2 AND B3) OR (NOT B0 AND B1 AND NOT B2);
    F <= (NOT B0 AND B2 AND B3) OR (NOT B0 AND NOT B1 AND B3) OR (NOT B0 AND NOT B1 AND B2) OR (B0 AND B1 AND NOT B2 AND B3);
    G <= (NOT B0 AND NOT B1 AND NOT B2) OR (NOT B0 AND B1 AND B2 AND B3) OR (B0 AND B1 AND NOT B2 AND NOT B3);
end Comportamento;